`timescale 1ns / 1ps

module decode_enb_leds(
    input [2:0] sel,
    output reg [7:0] enb_leds
    );

//
// Complete this block
//
endmodule
