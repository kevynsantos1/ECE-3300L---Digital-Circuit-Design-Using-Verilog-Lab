
module mult4 (
	     input [3:0] A, B,
	     output [7:0] X
	     );

//
// fill in the verilog code here to implement a 4-bit multiplier, 
// using multiple instances of the add4 module.
//   
   
endmodule // mult4

